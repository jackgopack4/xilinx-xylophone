module bus_interface_tb();

endmodule